library ieee;
use ieee.std_logic_1164.all;

entity INV_S_Box is

    port (a  : in  std_logic_vector(7 downto 0);
          temp : out std_logic_vector(7 downto 0));

end INV_S_Box;

architecture INV_S_Box_architecture of INV_S_Box is
Begin
 substitute: process(input) begin

        case a is

when x"00" => temp:= x"52";
when x"01" => temp := x"09";
when x"02" => temp:= x"6a";
when x"03" => temp := x"d5";
when x"04" => temp := x"30";
when x"05" => temp := x"36";
when x"06" => temp := x"a5";
when x"07" => temp := x"38";
when x"08" => temp := x"bf";
when x"09" => temp := x"40";
when x"0a" => temp := x"a3";
when x"0b" => temp := x"9e";
when x"0c" => temp := x"81";
when x"0d" => temp := x"f3";
when x"0e" => temp := x"d7";
when x"0f" => temp := x"fb";
when x"10" => temp := x"7c";
when x"11" => temp := x"e3";
when x"12" => temp := x"39";
when x"13" => temp := x"82";
when x"14" => temp := x"9b";
when x"15" => temp := x"2f";
when x"16" => temp := x"ff";
when x"17" => temp := x"87";
when x"18" => temp := x"34";
when x"19" => temp := x"8e";
when x"1a" => temp := x"43";
when x"1b" => temp := x"44";
when x"1c" => temp := x"c4";
when x"1d" => temp := x"de";
when x"1e" => temp := x"e9";
when x"1f" => temp := x"cb";
when x"20" => temp := x"54";
when x"21" => temp := x"7b";
when x"22" => temp := x"94";
when x"23" => temp := x"32";
when x"24" => temp := x"a6";
when x"25" => temp := x"c2";
when x"26" => temp := x"23";
when x"27" => temp := x"3d";
when x"28" => temp := x"ee";
when x"29" => temp := x"4c";
when x"2a" => temp := x"95";
when x"2b" => temp := x"0b";
when x"2c" => temp := x"42";
when x"2d" => temp := x"fa";
when x"2e" => temp := x"c3";
when x"2f" => temp := x"49";
when x"30" => temp := x"08";
when x"31" => temp := x"2e";
when x"32" => temp := x"a1";
when x"33" => temp := x"66";
when x"34" => temp := x"28";
when x"35" => temp := x"d9";
when x"36" => temp := x"24";
when x"37" => temp := x"b2";
when x"38" => temp := x"76";
when x"39" => temp := x"5b";
when x"3a" => temp := x"a2";
when x"3b" => temp := x"49";
when x"3c" => temp := x"6d";
when x"3d" => temp := x"8b";
when x"3e" => temp := x"d1";
when x"40" => temp := x"72";
when x"41" => temp := x"f8";
when x"42" => temp := x"f6";
when x"43" => temp := x"64";
when x"44" => temp := x"86";
when x"45" => temp := x"68";
when x"46" => temp := x"98";
when x"47" => temp := x"16";
when x"48" => temp := x"d4";
when x"49" => temp := x"a4";
when x"4a" => temp := x"5c";
when x"4b" => temp := x"cc";
when x"4c" => temp := x"5d";
when x"4d" => temp := x"65";
when x"4e" => temp := x"b6";
when x"4f" => temp := x"92";
when x"50" => temp := x"6c";
when x"51" => temp := x"70";
when x"52" => temp := x"48";
when x"53" => temp := x"50";
when x"54" => temp := x"fd";
when x"55" => temp := x"ed";
when x"56" => temp := x"b9";
when x"57" => temp := x"da";
when x"58" => temp := x"5e";
when x"59" => temp := x"15";
when x"5a" => temp := x"46";
when x"5b" => temp := x"57";
when x"5c" => temp := x"a7";
when x"5d" => temp := x"8d";
when x"5e" => temp := x"9d";
when x"5f" => temp := x"84";
when x"60" => temp := x"90";
when x"61" => temp := x"d8";
when x"62" => temp := x"ab";
when x"63" => temp := x"00";
when x"64" => temp := x"8c";
when x"65" => temp := x"bc";
when x"66" => temp := x"d3";
when x"67" => temp := x"0a";
when x"68" => temp := x"f7";
when x"69" => temp := x"e4";
when x"6a" => temp := x"58";
when x"6b" => temp := x"05";
when x"6c" => temp := x"b8";
when x"6d" => temp := x"b3";
when x"6e" => temp := x"45";
when x"6f" => temp := x"06";
when x"70" => temp := x"d0";
when x"71" => temp := x"2c";
when x"72" => temp := x"1e";
when x"73" => temp := x"8f";
when x"74" => temp := x"ca";
when x"75" => temp := x"3f";
when x"76" => temp := x"0f";
when x"77" => temp := x"02";
when x"78" => temp := x"c1";
when x"79" => temp := x"af";
when x"7a" => temp := x"bd";
when x"7b" => temp := x"03";
when x"7c" => temp := x"01";
when x"7d" => temp := x"13";
when x"7e" => temp := x"8a";
when x"7f" => temp := x"6b";
when x"80" => temp := x"3a";
when x"81" => temp := x"91";
when x"82" => temp := x"11";
when x"83" => temp := x"41";
when x"84" => temp := x"4f";
when x"85" => temp := x"67";
when x"86" => temp := x"dc";
when x"87" => temp := x"ea";
when x"88" => temp := x"97";
when x"89" => temp := x"f2";
when x"8a" => temp := x"cf";
when x"8b" => temp := x"ce";
when x"8c" => temp := x"f0";
when x"8d" => temp := x"b4";
when x"8e" => temp := x"e6";
when x"8f" => temp := x"73";
when x"90" => temp := x"96";
when x"91" => temp := x"ac";
when x"92" => temp := x"74";
when x"93" => temp := x"22";
when x"94" => temp := x"e7";
when x"95" => temp := x"ad";
when x"96" => temp := x"35";
when x"97" => temp := x"85";
when x"98" => temp := x"e2";
when x"99" => temp := x"f9";
when x"9a" => temp := x"37";
when x"9b" => temp := x"e8";
when x"9c" => temp := x"1c";
when x"9d" => temp := x"75";
when x"9e" => temp := x"df";
when x"9f" => temp := x"6e";
when x"a0" => temp := x"47";
when x"a1" => temp := x"f1";
when x"a2" => temp := x"1a";
when x"a3" => temp := x"71";
when x"a4" => temp := x"1d";
when x"a5" => temp := x"29";
when x"a6" => temp := x"c5";
when x"a7" => temp := x"89";
when x"a8" => temp := x"6f";
when x"a9" => temp := x"b7";
when x"aa" => temp := x"62";
when x"ab" => temp := x"0e";
when x"ac" => temp := x"aa";
when x"ad" => temp := x"18";
when x"ae" => temp := x"be";
when x"af" => temp := x"1b";
when x"b0" => temp := x"fc";
when x"b1" => temp := x"56";
when x"b2" => temp := x"3e";
when x"b3" => temp := x"4b";
when x"b4" => temp := x"c6";
when x"b5" => temp := x"d2";
when x"b6" => temp := x"79";
when x"b7" => temp := x"20";
when x"b8" => temp := x"9a";
when x"b9" => temp := x"db";
when x"ba" => temp := x"c0";
when x"bb" => temp := x"fe";
when x"bc" => temp := x"78";
when x"bd" => temp := x"cd";
when x"be" => temp := x"5a";
when x"bf" => temp := x"f4";
when x"c0" => temp := x"1f";
when x"c1" => temp := x"dd";
when x"c2" => temp := x"a8";
when x"c3" => temp := x"33";
when x"c4" => temp := x"88";
when x"c5" => temp := x"07";
when x"c6" => temp := x"c7";
when x"c7" => temp := x"31";
when x"c8" => temp := x"b1";
when x"c9" => temp := x"12";
when x"ca" => temp := x"10";
when x"cb" => temp := x"59";
when x"cc" => temp := x"27";
when x"cd" => temp := x"80";
when x"ce" => temp := x"ec";
when x"cf" => temp := x"5f";
when x"d0" => temp := x"60";
when x"d1" => temp := x"51";
when x"d2" => temp := x"7f";
when x"d3" => temp := x"a9";
when x"d4" => temp := x"19";
when x"d5" => temp := x"b5";
when x"d6" => temp := x"4a";
when x"d7" => temp := x"0d";
when x"d8" => temp := x"2d";
when x"d9" => temp := x"e5";
when x"da" => temp := x"7a";
when x"db" => temp := x"9f";
when x"dc" => temp := x"93";
when x"dd" => temp := x"c9";
when x"de" => temp := x"9c";
when x"df" => temp := x"ef";
when x"e0" => temp := x"a0";
when x"e1" => temp := x"e0";
when x"e2" => temp := x"3b";
when x"e3" => temp := x"4d";
when x"e4" => temp := x"ae";
when x"e5" => temp := x"2a";
when x"e6" => temp := x"f5";
when x"e7" => temp := x"b0";
when x"e8" => temp := x"c8";
when x"e9" => temp := x"eb";
when x"ea" => temp := x"bb";
when x"eb" => temp := x"3c";
when x"ec" => temp := x"83";
when x"ed" => temp := x"53";
when x"ee" => temp := x"99";
when x"ef" => temp := x"61";
when x"f0" => temp := x"17";
when x"f1" => temp := x"2b";
when x"f2" => temp := x"04";
when x"f3" => temp := x"7e";
when x"f4" => temp := x"ba";
when x"f5" => temp := x"77";
when x"f6" => temp := x"d6";
when x"f7" => temp := x"26";
when x"f8" => temp := x"e1";
when x"f9" => temp := x"69";
when x"fa" => temp := x"14";
when x"fb" => temp := x"63";
when x"fc" => temp := x"55";
when x"fd" => temp := x"21";
when x"fe" => temp := x"0c";
when x"ff" => temp := x"7d";
       when others => null;

        end case;

    end process;

end INV_S_Box_architecture;
